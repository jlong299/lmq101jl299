
module cnst_rom (
	address,
	clock,
	q);	

	input		address;
	input		clock;
	output	[7:0]	q;
endmodule
